localparam IDLE = 3'b000;
localparam CHECK_LEN = 3'b001;
localparam STREAM_IN = 3'b010;
localparam FIR_COMP = 3'b011;
localparam STREAM_OUT = 3'b100;
localparam DONE = 3'b101;
